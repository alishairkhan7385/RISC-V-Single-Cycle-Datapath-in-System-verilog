module control(cntrl_bits,breq,brlt,pc_sel,imm_sel,reg_wen,brUn,b_sel,a_sel,alu_sel,memRw,wb_sel,sw_imm_sel,lw_imm_sel);
input logic [8:0] cntrl_bits;
input logic breq;
input logic brlt;

output logic pc_sel; 
output logic [2:0] imm_sel;
output logic reg_wen;
output logic brUn;
output logic b_sel;
output logic a_sel;
output logic [3:0] alu_sel;
output logic memRw;
output logic [1:0] wb_sel;
output logic [1:0] sw_imm_sel;//sh,sb
output logic [2:0] lw_imm_sel;//lh,lb
always_comb
begin
	casez(cntrl_bits)
		9'b000001100://add
			begin
				pc_sel=1'b0;
				imm_sel=3'bxxx;
				reg_wen=1'b1;
				brUn=1'b0;
				b_sel=1'b0;
				a_sel=1'b0;
				alu_sel=4'b0000;
				memRw=1'b0;
				wb_sel=2'b01;
			end
			
		9'b100001100://sub
			begin
				pc_sel=1'b0;
				imm_sel=3'bxxx;
				reg_wen=1'b1;
				brUn=1'b0;
				b_sel=1'b0;
				a_sel=1'b0;
				alu_sel=4'b0010;
				memRw=1'b0;
				wb_sel=2'b01;
			end
			
		9'b010001100://xor
			begin
				pc_sel=1'b0;
				imm_sel=3'bxxx;
				reg_wen=1'b1;
				brUn=1'b0;
				b_sel=1'b0;
				a_sel=1'b0;
				alu_sel=4'b0011;
				memRw=1'b0;
				wb_sel=2'b01;
			end
			
		9'b011001100://or
			begin
				pc_sel=1'b0;
				imm_sel=3'bxxx;
				reg_wen=1'b1;
				brUn=1'b0;
				b_sel=1'b0;
				a_sel=1'b0;
				alu_sel=4'b0100;
				memRw=1'b0;
				wb_sel=2'b01;
			end
			
		9'b011101100://and
			begin
				pc_sel=1'b0;
				imm_sel=3'bxxx;
				reg_wen=1'b1;
				brUn=1'b0;
				b_sel=1'b0;
				a_sel=1'b0;
				alu_sel=4'b0101;
				memRw=1'b0;
				wb_sel=2'b01;
			end
		9'b000101100://sll
			begin
				pc_sel=1'b0;
				imm_sel=3'bxxx;
				reg_wen=1'b1;
				brUn=1'b0;
				b_sel=1'b0;
				a_sel=1'b0;
				alu_sel=4'b0110;
				memRw=1'b0;
				wb_sel=2'b01;
			end
		9'b010101100://srl
			begin
				pc_sel=1'b0;
				imm_sel=3'bxxx;
				reg_wen=1'b1;
				brUn=1'b0;
				b_sel=1'b0;
				a_sel=1'b0;
				alu_sel=4'b0111;
				memRw=1'b0;
				wb_sel=2'b01;
			end
		9'b110101100://sra
			begin
				pc_sel=1'b0;
				imm_sel=3'bxxx;
				reg_wen=1'b1;
				brUn=1'b0;
				b_sel=1'b0;
				a_sel=1'b0;
				alu_sel=4'b1000;
				memRw=1'b0;
				wb_sel=2'b01;
			end
		
		9'b001001100://slt
			begin
				pc_sel=1'b0;
				imm_sel=3'bxxx;
				reg_wen=1'b1;
				brUn=1'b0;
				b_sel=1'b0;
				a_sel=1'b0;
				alu_sel=4'b1001;
				memRw=1'b0;
				wb_sel=2'b01;
			end
		9'b001101100://sltu
			begin
				pc_sel=1'b0;
				imm_sel=3'bxxx;
				reg_wen=1'b1;
				brUn=1'b0;
				b_sel=1'b0;
				a_sel=1'b0;
				alu_sel=4'b1010;
				memRw=1'b0;
				wb_sel=2'b01;
			end
		//I type
		9'bz00000100://addi
			begin
				pc_sel=1'b0;
				imm_sel=3'b000;
				reg_wen=1'b1;
				brUn=1'b0;
				b_sel=1'b1;
				a_sel=1'b0;
				alu_sel=4'b0000;
				memRw=1'b0;
				wb_sel=2'b01;
			end
		
		9'bz100000100://xori
			begin
				pc_sel=1'b0;
				imm_sel=3'b000;
				reg_wen=1'b1;
				brUn=1'b0;
				b_sel=1'b1;
				a_sel=1'b0;
				alu_sel=4'b0011;
				memRw=1'b0;
				wb_sel=2'b01;
			end
		
		9'bz110000100://ori
			begin
				pc_sel=1'b0;
				imm_sel=3'b000;
				reg_wen=1'b1;
				brUn=1'b0;
				b_sel=1'b1;
				a_sel=1'b0;
				alu_sel=4'b0100;
				memRw=1'b0;
				wb_sel=2'b01;
			end
		
		9'bz11100100://andi
			begin
				pc_sel=1'b0;
				imm_sel=3'b000;
				reg_wen=1'b1;
				brUn=1'b0;
				b_sel=1'b1;
				a_sel=1'b0;
				alu_sel=4'b0101;
				memRw=1'b0;
				wb_sel=2'b01;
			end
		9'bz01000100://slti
			begin
				pc_sel=1'b0;
				imm_sel=3'b000;
				reg_wen=1'b1;
				brUn=1'b0;
				b_sel=1'b1;
				a_sel=1'b0;
				alu_sel=4'b1001;
				memRw=1'b0;
				wb_sel=2'b01;
			end
		9'bz01100100://sltiu
			begin
				pc_sel=1'b0;
				imm_sel=3'b000;
				reg_wen=1'b1;
				brUn=1'b0;
				b_sel=1'b1;
				a_sel=1'b0;
				alu_sel=4'b1010;
				memRw=1'b0;
				wb_sel=2'b01;
			end
		9'bz10000100://xori
			begin
				pc_sel=1'b0;
				imm_sel=3'b000;
				reg_wen=1'b1;
				brUn=1'b0;
				b_sel=1'b1;
				a_sel=1'b0;
				alu_sel=4'b0011;
				memRw=1'b0;
				wb_sel=2'b01;
			end
		9'bz11000100://ori
			begin
				pc_sel=1'b0;
				imm_sel=3'b000;
				reg_wen=1'b1;
				brUn=1'b0;
				b_sel=1'b1;
				a_sel=1'b0;
				alu_sel=4'b0100;
				memRw=1'b0;
				wb_sel=2'b01;
			end
		9'b000100100://slli
			begin
				pc_sel=1'b0;
				imm_sel=3'b101;
				reg_wen=1'b1;
				brUn=1'b0;
				b_sel=1'b1;
				a_sel=1'b0;
				alu_sel=4'b0110;
				memRw=1'b0;
				wb_sel=2'b01;
			end
		9'b010100100://srli
			begin
				pc_sel=1'b0;
				imm_sel=3'b101;
				reg_wen=1'b1;
				brUn=1'b0;
				b_sel=1'b1;
				a_sel=1'b0;
				alu_sel=4'b0111;
				memRw=1'b0;
				wb_sel=2'b01;
			end
		9'b110100100://srai
			begin
				pc_sel=1'b0;
				imm_sel=3'b101;
				reg_wen=1'b1;
				brUn=1'b0;
				b_sel=1'b1;
				a_sel=1'b0;
				alu_sel=4'b1000;
				memRw=1'b0;
				wb_sel=2'b01;
			end
			
		9'bz01001000://sw
			begin
				pc_sel=1'b0;
				imm_sel=3'b001;
				reg_wen=1'b0;
				brUn=1'b0;
				b_sel=1'b1;
				a_sel=1'b0;
				alu_sel=4'b0000;
				memRw=1'b1;
				wb_sel=2'bxx;
				sw_imm_sel=2'b00;
			end
		9'bz00001000://sb
			begin
				pc_sel=1'b0;
				imm_sel=3'b001;
				reg_wen=1'b0;
				brUn=1'b0;
				b_sel=1'b1;
				a_sel=1'b0;
				alu_sel=4'b0000;
				memRw=1'b1;
				wb_sel=2'bxx;
				sw_imm_sel=2'b01;
			end
		9'bz00101000://sh
			begin
				pc_sel=1'b0;
				imm_sel=3'b001;
				reg_wen=1'b0;
				brUn=1'b0;
				b_sel=1'b1;
				a_sel=1'b0;
				alu_sel=4'b0000;
				memRw=1'b1;
				sw_imm_sel=2'b10;
			end
		9'bz01000000://lw
			begin
				pc_sel=1'b0;
				imm_sel=3'b000;
				reg_wen=1'b1;
				brUn=1'b0;
				b_sel=1'b1;
				a_sel=1'b0;
				alu_sel=4'b0000;
				memRw=1'b0;
				wb_sel=2'b00;
				lw_imm_sel=3'b000;
			end
		9'bz00100000://lh
			begin
				pc_sel=1'b0;
				imm_sel=3'b000;
				reg_wen=1'b1;
				brUn=1'b0;
				b_sel=1'b1;
				a_sel=1'b0;
				alu_sel=4'b0000;
				memRw=1'b0;
				wb_sel=2'b00;
				lw_imm_sel=3'b001;
			end
		9'bz00000000://lb
			begin
				pc_sel=1'b0;
				imm_sel=3'b000;
				reg_wen=1'b1;
				brUn=1'b0;
				b_sel=1'b1;
				a_sel=1'b0;
				alu_sel=4'b0000;
				memRw=1'b0;
				wb_sel=2'b00;
				lw_imm_sel=3'b010;
			end
		9'bz10100000://lhu
			begin
				pc_sel=1'b0;
				imm_sel=3'b000;
				reg_wen=1'b1;
				brUn=1'b0;
				b_sel=1'b1;
				a_sel=1'b0;
				alu_sel=4'b0000;
				memRw=1'b0;
				wb_sel=2'b00;
				lw_imm_sel=3'b011;
			end
		9'bz10000000://lbu
			begin
				pc_sel=1'b0;
				imm_sel=3'b000;
				reg_wen=1'b1;
				brUn=1'b0;
				b_sel=1'b1;
				a_sel=1'b0;
				alu_sel=4'b0000;
				memRw=1'b0;
				wb_sel=2'b00;
				lw_imm_sel=3'b100;
			end
		//branch
		9'bz00011000://beq
			begin
				pc_sel=breq?1:0;
				imm_sel=3'b010;
				reg_wen=1'b0;
				brUn=1'b0;
				b_sel=1'b1;
				a_sel=1'b1;
				alu_sel=4'b0000;
				memRw=1'b0;
				wb_sel=2'bxx;
			end
		9'bz00111000://bne
			begin
				pc_sel=breq?0:1;
				imm_sel=3'b010;
				reg_wen=1'b0;
				brUn=1'b0;
				b_sel=1'b1;
				a_sel=1'b1;
				alu_sel=4'b0000;
				memRw=1'b0;
				wb_sel=2'bxx;
			end
		9'bz10011000://blt
			begin
				pc_sel=brlt?1:0;
				imm_sel=3'b010;
				reg_wen=1'b0;
				brUn=1'b0;
				b_sel=1'b1;
				a_sel=1'b1;
				alu_sel=4'b0000;
				memRw=1'b0;
				wb_sel=2'bxx;
			end
		9'bz10111000://bge
			begin
				pc_sel=(breq||~brlt)?1:0;
				imm_sel=3'b010;
				reg_wen=1'b0;
				brUn=1'b0;
				b_sel=1'b1;
				a_sel=1'b1;
				alu_sel=4'b0000;
				memRw=1'b0;
				wb_sel=2'bxx;
			end
		9'bz11011000://bltu
			begin
				pc_sel=brlt?1:0;
				imm_sel=3'b010;
				reg_wen=1'b0;
				brUn=1'b1;
				b_sel=1'b1;
				a_sel=1'b1;
				alu_sel=4'b0000;
				memRw=1'b0;
				wb_sel=2'bxx;
			end
		9'bz11111000://bgeu
			begin
				pc_sel=(breq||~brlt)?1:0;
				imm_sel=3'b010;
				reg_wen=1'b0;
				brUn=1'b1;
				b_sel=1'b1;
				a_sel=1'b1;
				alu_sel=4'b0000;
				memRw=1'b0;
				wb_sel=2'bxx;
			end
		9'bzzzz11011://jal
			begin
				pc_sel=1'b1;
				imm_sel=3'b011;
				reg_wen=1'b1;
				brUn=1'b0;
				b_sel=1'b1;
				a_sel=1'b1;
				alu_sel=4'b0000;
				memRw=1'b0;
				wb_sel=2'b10;
			end
		9'bz00011001://jalr
			begin
				pc_sel=1'b1;
				imm_sel=3'b000;
				reg_wen=1'b1;
				brUn=1'b0;
				b_sel=1'b1;
				a_sel=1'b0;
				alu_sel=4'b0000;
				memRw=1'b0;
				wb_sel=2'b10;
			end	
		9'bzzzz01101://lui
			begin
				pc_sel=1'b0;
				imm_sel=3'b100;
				reg_wen=1'b1;
				brUn=1'bx;
				b_sel=1'b0;
				a_sel=1'b0;
				alu_sel=4'b0000;
				memRw=1'b0;
				wb_sel=2'b11;
			end
		9'bzzzz00101://auipc
			begin
				pc_sel=1'b0;
				imm_sel=3'b100;
				reg_wen=1'b1;
				brUn=1'bx;
				b_sel=1'b1;
				a_sel=1'b1;
				alu_sel=4'b0000;
				memRw=1'b0;
				wb_sel=2'b01;
			end
	endcase
end
endmodule
